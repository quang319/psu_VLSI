module widthCb (
	input wire [7:0] Y,

	output reg [31:0] result
	);

	always @(Y) begin
		case (Y)
			8'd0: result = 32'h0004ded0; 
			8'd1: result = 32'h0004ece3; 
			8'd2: result = 32'h0004faf6; 
			8'd3: result = 32'h00050909; 
			8'd4: result = 32'h0005171c; 
			8'd5: result = 32'h0005252f; 
			8'd6: result = 32'h00053342; 
			8'd7: result = 32'h00054155; 
			8'd8: result = 32'h00054f68; 
			8'd9: result = 32'h00055d7b; 
			8'd10: result = 32'h00056b8e; 
			8'd11: result = 32'h000579a1; 
			8'd12: result = 32'h000587b4; 
			8'd13: result = 32'h000595c7; 
			8'd14: result = 32'h0005a3da; 
			8'd15: result = 32'h0005b1ed; 
			8'd16: result = 32'h0005c000; 
			8'd17: result = 32'h0005ce12; 
			8'd18: result = 32'h0005dc25; 
			8'd19: result = 32'h0005ea38; 
			8'd20: result = 32'h0005f84b; 
			8'd21: result = 32'h0006065e; 
			8'd22: result = 32'h00061471; 
			8'd23: result = 32'h00062284; 
			8'd24: result = 32'h00063097; 
			8'd25: result = 32'h00063eaa; 
			8'd26: result = 32'h00064cbd; 
			8'd27: result = 32'h00065ad0; 
			8'd28: result = 32'h000668e3; 
			8'd29: result = 32'h000676f6; 
			8'd30: result = 32'h00068509; 
			8'd31: result = 32'h0006931c; 
			8'd32: result = 32'h0006a12f; 
			8'd33: result = 32'h0006af42; 
			8'd34: result = 32'h0006bd55; 
			8'd35: result = 32'h0006cb68; 
			8'd36: result = 32'h0006d97b; 
			8'd37: result = 32'h0006e78e; 
			8'd38: result = 32'h0006f5a1; 
			8'd39: result = 32'h000703b4; 
			8'd40: result = 32'h000711c7; 
			8'd41: result = 32'h00071fda; 
			8'd42: result = 32'h00072ded; 
			8'd43: result = 32'h00073c00; 
			8'd44: result = 32'h00074a13; 
			8'd45: result = 32'h00075826; 
			8'd46: result = 32'h00076639; 
			8'd47: result = 32'h0007744c; 
			8'd48: result = 32'h0007825f; 
			8'd49: result = 32'h00079072; 
			8'd50: result = 32'h00079e85; 
			8'd51: result = 32'h0007ac98; 
			8'd52: result = 32'h0007baab; 
			8'd53: result = 32'h0007c8be; 
			8'd54: result = 32'h0007d6d1; 
			8'd55: result = 32'h0007e4e4; 
			8'd56: result = 32'h0007f2f7; 
			8'd57: result = 32'h0008010a; 
			8'd58: result = 32'h00080f1d; 
			8'd59: result = 32'h00081d30; 
			8'd60: result = 32'h00082b42; 
			8'd61: result = 32'h00083955; 
			8'd62: result = 32'h00084768; 
			8'd63: result = 32'h0008557b; 
			8'd64: result = 32'h0008638e; 
			8'd65: result = 32'h000871a1; 
			8'd66: result = 32'h00087fb4; 
			8'd67: result = 32'h00088dc7; 
			8'd68: result = 32'h00089bda; 
			8'd69: result = 32'h0008a9ed; 
			8'd70: result = 32'h0008b800; 
			8'd71: result = 32'h0008c613; 
			8'd72: result = 32'h0008d426; 
			8'd73: result = 32'h0008e239; 
			8'd74: result = 32'h0008f04c; 
			8'd75: result = 32'h0008fe5f; 
			8'd76: result = 32'h00090c72; 
			8'd77: result = 32'h00091a85; 
			8'd78: result = 32'h00092898; 
			8'd79: result = 32'h000936ab; 
			8'd80: result = 32'h000944be; 
			8'd81: result = 32'h000952d1; 
			8'd82: result = 32'h000960e4; 
			8'd83: result = 32'h00096ef7; 
			8'd84: result = 32'h00097d0a; 
			8'd85: result = 32'h00098b1d; 
			8'd86: result = 32'h00099930; 
			8'd87: result = 32'h0009a743; 
			8'd88: result = 32'h0009b556; 
			8'd89: result = 32'h0009c369; 
			8'd90: result = 32'h0009d17c; 
			8'd91: result = 32'h0009df8f; 
			8'd92: result = 32'h0009eda2; 
			8'd93: result = 32'h0009fbb5; 
			8'd94: result = 32'h000a09c8; 
			8'd95: result = 32'h000a17db; 
			8'd96: result = 32'h000a25ee; 
			8'd97: result = 32'h000a3401; 
			8'd98: result = 32'h000a4214; 
			8'd99: result = 32'h000a5027; 
			8'd100: result = 32'h000a5e3a; 
			8'd101: result = 32'h000a6c4d; 
			8'd102: result = 32'h000a7a60; 
			8'd103: result = 32'h000a8872; 
			8'd104: result = 32'h000a9685; 
			8'd105: result = 32'h000aa498; 
			8'd106: result = 32'h000ab2ab; 
			8'd107: result = 32'h000ac0be; 
			8'd108: result = 32'h000aced1; 
			8'd109: result = 32'h000adce4; 
			8'd110: result = 32'h000aeaf7; 
			8'd111: result = 32'h000af90a; 
			8'd112: result = 32'h000b071d; 
			8'd113: result = 32'h000b1530; 
			8'd114: result = 32'h000b2343; 
			8'd115: result = 32'h000b3156; 
			8'd116: result = 32'h000b3f69; 
			8'd117: result = 32'h000b4d7c; 
			8'd118: result = 32'h000b5b8f; 
			8'd119: result = 32'h000b69a2; 
			8'd120: result = 32'h000b77b5; 
			8'd121: result = 32'h000b85c8; 
			8'd122: result = 32'h000b93db; 
			8'd123: result = 32'h000ba1ee; 
			8'd124: result = 32'h000bb001; 
			8'd125: result = 32'h000bbe14; 
			8'd126: result = 32'h00000000; 
			8'd127: result = 32'h00000000; 
			8'd128: result = 32'h00000000; 
			8'd129: result = 32'h00000000; 
			8'd130: result = 32'h00000000; 
			8'd131: result = 32'h00000000; 
			8'd132: result = 32'h00000000; 
			8'd133: result = 32'h00000000; 
			8'd134: result = 32'h00000000; 
			8'd135: result = 32'h00000000; 
			8'd136: result = 32'h00000000; 
			8'd137: result = 32'h00000000; 
			8'd138: result = 32'h00000000; 
			8'd139: result = 32'h00000000; 
			8'd140: result = 32'h00000000; 
			8'd141: result = 32'h00000000; 
			8'd142: result = 32'h00000000; 
			8'd143: result = 32'h00000000; 
			8'd144: result = 32'h00000000; 
			8'd145: result = 32'h00000000; 
			8'd146: result = 32'h00000000; 
			8'd147: result = 32'h00000000; 
			8'd148: result = 32'h00000000; 
			8'd149: result = 32'h00000000; 
			8'd150: result = 32'h00000000; 
			8'd151: result = 32'h00000000; 
			8'd152: result = 32'h00000000; 
			8'd153: result = 32'h00000000; 
			8'd154: result = 32'h00000000; 
			8'd155: result = 32'h00000000; 
			8'd156: result = 32'h00000000; 
			8'd157: result = 32'h00000000; 
			8'd158: result = 32'h00000000; 
			8'd159: result = 32'h00000000; 
			8'd160: result = 32'h00000000; 
			8'd161: result = 32'h00000000; 
			8'd162: result = 32'h00000000; 
			8'd163: result = 32'h00000000; 
			8'd164: result = 32'h00000000; 
			8'd165: result = 32'h00000000; 
			8'd166: result = 32'h00000000; 
			8'd167: result = 32'h00000000; 
			8'd168: result = 32'h00000000; 
			8'd169: result = 32'h00000000; 
			8'd170: result = 32'h00000000; 
			8'd171: result = 32'h00000000; 
			8'd172: result = 32'h00000000; 
			8'd173: result = 32'h00000000; 
			8'd174: result = 32'h00000000; 
			8'd175: result = 32'h00000000; 
			8'd176: result = 32'h00000000; 
			8'd177: result = 32'h00000000; 
			8'd178: result = 32'h00000000; 
			8'd179: result = 32'h00000000; 
			8'd180: result = 32'h00000000; 
			8'd181: result = 32'h00000000; 
			8'd182: result = 32'h00000000; 
			8'd183: result = 32'h00000000; 
			8'd184: result = 32'h00000000; 
			8'd185: result = 32'h00000000; 
			8'd186: result = 32'h00000000; 
			8'd187: result = 32'h00000000; 
			8'd188: result = 32'h000bbe14; 
			8'd189: result = 32'h000b912f; 
			8'd190: result = 32'h000b644a; 
			8'd191: result = 32'h000b3764; 
			8'd192: result = 32'h000b0a7f; 
			8'd193: result = 32'h000add9a; 
			8'd194: result = 32'h000ab0b5; 
			8'd195: result = 32'h000a83d0; 
			8'd196: result = 32'h000a56ea; 
			8'd197: result = 32'h000a2a05; 
			8'd198: result = 32'h0009fd20; 
			8'd199: result = 32'h0009d03b; 
			8'd200: result = 32'h0009a356; 
			8'd201: result = 32'h00097670; 
			8'd202: result = 32'h0009498b; 
			8'd203: result = 32'h00091ca6; 
			8'd204: result = 32'h0008efc1; 
			8'd205: result = 32'h0008c2dc; 
			8'd206: result = 32'h000895f6; 
			8'd207: result = 32'h00086911; 
			8'd208: result = 32'h00083c2c; 
			8'd209: result = 32'h00080f47; 
			8'd210: result = 32'h0007e262; 
			8'd211: result = 32'h0007b57c; 
			8'd212: result = 32'h00078897; 
			8'd213: result = 32'h00075bb2; 
			8'd214: result = 32'h00072ecd; 
			8'd215: result = 32'h000701e8; 
			8'd216: result = 32'h0006d502; 
			8'd217: result = 32'h0006a81d; 
			8'd218: result = 32'h00067b38; 
			8'd219: result = 32'h00064e53; 
			8'd220: result = 32'h0006216e; 
			8'd221: result = 32'h0005f488; 
			8'd222: result = 32'h0005c7a3; 
			8'd223: result = 32'h00059abe; 
			8'd224: result = 32'h00056dd9; 
			8'd225: result = 32'h000540f4; 
			8'd226: result = 32'h0005140e; 
			8'd227: result = 32'h0004e729; 
			8'd228: result = 32'h0004ba44; 
			8'd229: result = 32'h00048d5f; 
			8'd230: result = 32'h0004607a; 
			8'd231: result = 32'h00043394; 
			8'd232: result = 32'h000406af; 
			8'd233: result = 32'h0003d9ca; 
			8'd234: result = 32'h0003ace5; 
			8'd235: result = 32'h00038000; 
			8'd236: result = 32'h0003531a; 
			8'd237: result = 32'h00032635; 
			8'd238: result = 32'h0002f950; 
			8'd239: result = 32'h0002cc6b; 
			8'd240: result = 32'h00029f85; 
			8'd241: result = 32'h000272a0; 
			8'd242: result = 32'h000245bb; 
			8'd243: result = 32'h000218d6; 
			8'd244: result = 32'h0001ebf1; 
			8'd245: result = 32'h0001bf0b; 
			8'd246: result = 32'h00019226; 
			8'd247: result = 32'h00016541; 
			8'd248: result = 32'h0001385c; 
			8'd249: result = 32'h00010b77; 
			8'd250: result = 32'h0000de91; 
			8'd251: result = 32'h0000b1ac; 
			8'd252: result = 32'h000084c7; 
			8'd253: result = 32'h000057e2; 
			8'd254: result = 32'h00002afd; 
			8'd255: result = 32'hfffffe18; 

			default : result = 32'h00000000;
		endcase
	end

endmodule