
`define SKINTONE_IMAGE_INFO_BASE_FLOWID_FIELD				9:0
`define SKINTONE_IMAGE_INFO_WIDTH_FIELD						21:10
`define SKINTONE_IMAGE_INFO_HEIGHT_FIELD					33:22
`define SKINTONE_IMAGE_INFO_TYPE_FIELD						39:34
`define SKINTONE_IMAGE_INFO_FORMAT_FIELD					47:40
`define SKINTONE_IMAGE_INFO_FORMAT_COLOR_FIELD				43:40
`define SKINTONE_IMAGE_INFO_FORMAT_DEPTH_FIELD				47:44
`define SKINTONE_IMAGE_INFO_ACCUM_DEVICE_ID_FIELD			63:48
`define SKINTONE_IMAGE_INFO_ACCUM_ADDRESS_FIELD				127:64

`define AIM_NOTIFICATION_TARGET_DEVICE_ID_FIELD				15:0
`define SKINTONE_DATAPATH_STATUS_PIXEL_QUEUE_COUNT			17:0
`define SKINTONE_DATAPATH_STATUS_OUTPUT_QUEUE_COUNT			35:18	
			
`define SKINTONE_TAG_INDEX_PIXEL_FETCH						0
`define SKINTONE_TAG_INDEX_RESULT_STORE 					1
`define SKINTONE_TAG_INDEX_CONTROLLER 						2

