`ifndef _projectHeader_vh_
`define _projectHeader_vh_

`define ECy 32'h00009a3d
`define WL_Cb 32'h0005c000
`define ECx 32'h00006666
`define InvA 32'h00000285
`define K_l 32'h001f4000
`define InvB 32'h0000048f
`define WH_Cb 32'h00038000
`define NSint 32'hffffdb41
`define W_Cr 32'h0009b0a3
`define Cost 32'hffffcb9a
`define Y_max 32'h003ac000
`define Y_min 32'h00040000
`define WH_Cr 32'h00028000
`define fac 32'h007f8000
`define Radius 32'h00002000
`define Sint 32'h000024bf
`define Cy 32'h00260147
`define W_Cb 32'h000bbe14
`define WL_Cr 32'h00050000
`define Cx 32'h001b5851
`define K_h 32'h002f0000

`endif //_projectHeader_vh_